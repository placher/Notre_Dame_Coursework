module top_display(
	input [3:0] s,
	output reg [6:0] f);
	
	always @(s) begin
		case (s)
			4'b0000: f = 7'b1000000;
			4'b0001: f = 7'b1111001;
			4'b0010: f = 7'b0100100;
			4'b0011: f = 7'b0110000;
			4'b0100: f = 7'b0011001;
			4'b0101: f = 7'b0010010;
			4'b0110: f = 7'b0000010;
			4'b0111: f = 7'b1111000;
			4'b1000: f = 7'b0000000;
			4'b1001: f = 7'b0011000;
			4'b1010: f = 7'b0001000;
			4'b1011: f = 7'b0000011;
			4'b1100: f = 7'b1000110;
			4'b1101: f = 7'b0100001;
			4'b1110: f = 7'b0000110;
			4'b1111: f = 7'b0001110;
		endcase
	end
	
endmodule