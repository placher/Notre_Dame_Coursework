`timescale 1 ns/1 ns

module full_adder_tb();
	reg a, b, cin;
	wire cout, s;
	
	full_adder uut(a, b, cin, cout, s);
	
	initial begin
			 a = 0; b = 0; cin = 0;
		#10 a = 0; b = 0; cin = 1;
		#10 a = 0; b = 1; cin = 0;
		#10 a = 0; b = 1; cin = 1;
		#10 a = 1; b = 0; cin = 0;
		#10 a = 1; b = 0; cin = 1;
		#10 a = 1; b = 1; cin = 0;
		#10 a = 1; b = 1; cin = 1;
		#10;
	end

endmodule